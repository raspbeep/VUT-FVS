package sv_timer_t_gm_pkg;
    import uvm_pkg::*;
    import sv_param_pkg::*;
    import sv_timer_t_agent_pkg::*;

    `include "uvm_macros.svh"
    `include "golden_model.svh"
endpackage: sv_timer_t_gm_pkg
