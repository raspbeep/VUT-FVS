package sv_timer_t_agent_pkg;
    import uvm_pkg::*;
    import sv_param_pkg::*;

    `include "uvm_macros.svh"
    `include "transaction.svh"
    `include "monitor.svh"
    `include "coverage.svh"
    `include "driver.svh"
    `include "sequencer.svh"
    `include "sequence.svh"
    `include "agent.svh"
endpackage: sv_timer_t_agent_pkg
