package sv_timer_t_env_pkg;
    import uvm_pkg::*;
    import sv_param_pkg::*;
    import sv_timer_t_agent_pkg::*;
    import sv_timer_t_gm_pkg::*;

    `include "uvm_macros.svh"
    `include "scoreboard.svh"
    `include "env.svh"
endpackage: sv_timer_t_env_pkg
