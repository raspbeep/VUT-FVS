package sv_timer_t_test_pkg;
    import uvm_pkg::*;
    import sv_param_pkg::*;
    import sv_timer_t_agent_pkg::*;
    import sv_timer_t_gm_pkg::*;
    import sv_timer_t_env_pkg::*;

    `include "uvm_macros.svh"
    `include "test_base.svh"
    `include "test.svh"
endpackage: sv_timer_t_test_pkg
